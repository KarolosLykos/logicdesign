library verilog;
use verilog.vl_types.all;
entity myand_test is
end myand_test;
