library verilog;
use verilog.vl_types.all;
entity decoder2_2_4_struct is
    port(
        s1              : in     vl_logic;
        s0              : in     vl_logic;
        o0              : out    vl_logic;
        o1              : out    vl_logic;
        o2              : out    vl_logic;
        o3              : out    vl_logic
    );
end decoder2_2_4_struct;
