library verilog;
use verilog.vl_types.all;
entity testhier is
end testhier;
