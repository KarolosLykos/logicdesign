library verilog;
use verilog.vl_types.all;
entity test_all_xor is
end test_all_xor;
