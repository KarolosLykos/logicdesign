library verilog;
use verilog.vl_types.all;
entity testham is
end testham;
