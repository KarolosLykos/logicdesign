library verilog;
use verilog.vl_types.all;
entity test_all_dec is
end test_all_dec;
