library verilog;
use verilog.vl_types.all;
entity circuit3_2_test is
end circuit3_2_test;
