library verilog;
use verilog.vl_types.all;
entity circuit3_1 is
    port(
        a               : in     vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        z               : out    vl_logic
    );
end circuit3_1;
