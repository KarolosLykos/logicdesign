library verilog;
use verilog.vl_types.all;
entity decoder_test is
end decoder_test;
