library verilog;
use verilog.vl_types.all;
entity circuit3_1_test is
end circuit3_1_test;
